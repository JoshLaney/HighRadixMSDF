module DUTtester()
   input clk,
	