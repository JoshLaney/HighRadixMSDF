// soc_system.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module soc_system (
		input  wire        clk_clk,                               //             clk.clk
		output wire        hps_0_h2f_reset_reset_n,               // hps_0_h2f_reset.reset_n
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CLK, //    hps_0_hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD0,   //                .hps_io_emac1_inst_TXD0
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD1,   //                .hps_io_emac1_inst_TXD1
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD2,   //                .hps_io_emac1_inst_TXD2
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD3,   //                .hps_io_emac1_inst_TXD3
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD0,   //                .hps_io_emac1_inst_RXD0
		inout  wire        hps_0_hps_io_hps_io_emac1_inst_MDIO,   //                .hps_io_emac1_inst_MDIO
		output wire        hps_0_hps_io_hps_io_emac1_inst_MDC,    //                .hps_io_emac1_inst_MDC
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CTL, //                .hps_io_emac1_inst_RX_CTL
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CTL, //                .hps_io_emac1_inst_TX_CTL
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CLK, //                .hps_io_emac1_inst_RX_CLK
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD1,   //                .hps_io_emac1_inst_RXD1
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD2,   //                .hps_io_emac1_inst_RXD2
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD3,   //                .hps_io_emac1_inst_RXD3
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO0,     //                .hps_io_qspi_inst_IO0
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO1,     //                .hps_io_qspi_inst_IO1
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO2,     //                .hps_io_qspi_inst_IO2
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO3,     //                .hps_io_qspi_inst_IO3
		output wire        hps_0_hps_io_hps_io_qspi_inst_SS0,     //                .hps_io_qspi_inst_SS0
		output wire        hps_0_hps_io_hps_io_qspi_inst_CLK,     //                .hps_io_qspi_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_CMD,     //                .hps_io_sdio_inst_CMD
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D0,      //                .hps_io_sdio_inst_D0
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D1,      //                .hps_io_sdio_inst_D1
		output wire        hps_0_hps_io_hps_io_sdio_inst_CLK,     //                .hps_io_sdio_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D2,      //                .hps_io_sdio_inst_D2
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D3,      //                .hps_io_sdio_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D0,      //                .hps_io_usb1_inst_D0
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D1,      //                .hps_io_usb1_inst_D1
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D2,      //                .hps_io_usb1_inst_D2
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D3,      //                .hps_io_usb1_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D4,      //                .hps_io_usb1_inst_D4
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D5,      //                .hps_io_usb1_inst_D5
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D6,      //                .hps_io_usb1_inst_D6
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D7,      //                .hps_io_usb1_inst_D7
		input  wire        hps_0_hps_io_hps_io_usb1_inst_CLK,     //                .hps_io_usb1_inst_CLK
		output wire        hps_0_hps_io_hps_io_usb1_inst_STP,     //                .hps_io_usb1_inst_STP
		input  wire        hps_0_hps_io_hps_io_usb1_inst_DIR,     //                .hps_io_usb1_inst_DIR
		input  wire        hps_0_hps_io_hps_io_usb1_inst_NXT,     //                .hps_io_usb1_inst_NXT
		output wire        hps_0_hps_io_hps_io_spim0_inst_CLK,    //                .hps_io_spim0_inst_CLK
		output wire        hps_0_hps_io_hps_io_spim0_inst_MOSI,   //                .hps_io_spim0_inst_MOSI
		input  wire        hps_0_hps_io_hps_io_spim0_inst_MISO,   //                .hps_io_spim0_inst_MISO
		output wire        hps_0_hps_io_hps_io_spim0_inst_SS0,    //                .hps_io_spim0_inst_SS0
		input  wire        hps_0_hps_io_hps_io_uart0_inst_RX,     //                .hps_io_uart0_inst_RX
		output wire        hps_0_hps_io_hps_io_uart0_inst_TX,     //                .hps_io_uart0_inst_TX
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SDA,     //                .hps_io_i2c0_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SCL,     //                .hps_io_i2c0_inst_SCL
		input  wire        hps_0_hps_io_hps_io_can0_inst_RX,      //                .hps_io_can0_inst_RX
		output wire        hps_0_hps_io_hps_io_can0_inst_TX,      //                .hps_io_can0_inst_TX
		output wire        hps_0_hps_io_hps_io_trace_inst_CLK,    //                .hps_io_trace_inst_CLK
		output wire        hps_0_hps_io_hps_io_trace_inst_D0,     //                .hps_io_trace_inst_D0
		output wire        hps_0_hps_io_hps_io_trace_inst_D1,     //                .hps_io_trace_inst_D1
		output wire        hps_0_hps_io_hps_io_trace_inst_D2,     //                .hps_io_trace_inst_D2
		output wire        hps_0_hps_io_hps_io_trace_inst_D3,     //                .hps_io_trace_inst_D3
		output wire        hps_0_hps_io_hps_io_trace_inst_D4,     //                .hps_io_trace_inst_D4
		output wire        hps_0_hps_io_hps_io_trace_inst_D5,     //                .hps_io_trace_inst_D5
		output wire        hps_0_hps_io_hps_io_trace_inst_D6,     //                .hps_io_trace_inst_D6
		output wire        hps_0_hps_io_hps_io_trace_inst_D7,     //                .hps_io_trace_inst_D7
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO09,  //                .hps_io_gpio_inst_GPIO09
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO35,  //                .hps_io_gpio_inst_GPIO35
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO41,  //                .hps_io_gpio_inst_GPIO41
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO42,  //                .hps_io_gpio_inst_GPIO42
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO43,  //                .hps_io_gpio_inst_GPIO43
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO44,  //                .hps_io_gpio_inst_GPIO44
		output wire [14:0] memory_mem_a,                          //          memory.mem_a
		output wire [2:0]  memory_mem_ba,                         //                .mem_ba
		output wire        memory_mem_ck,                         //                .mem_ck
		output wire        memory_mem_ck_n,                       //                .mem_ck_n
		output wire        memory_mem_cke,                        //                .mem_cke
		output wire        memory_mem_cs_n,                       //                .mem_cs_n
		output wire        memory_mem_ras_n,                      //                .mem_ras_n
		output wire        memory_mem_cas_n,                      //                .mem_cas_n
		output wire        memory_mem_we_n,                       //                .mem_we_n
		output wire        memory_mem_reset_n,                    //                .mem_reset_n
		inout  wire [39:0] memory_mem_dq,                         //                .mem_dq
		inout  wire [4:0]  memory_mem_dqs,                        //                .mem_dqs
		inout  wire [4:0]  memory_mem_dqs_n,                      //                .mem_dqs_n
		output wire        memory_mem_odt,                        //                .mem_odt
		output wire [4:0]  memory_mem_dm,                         //                .mem_dm
		input  wire        memory_oct_rzqin,                      //                .oct_rzqin
		input  wire        reset_reset_n                          //           reset.reset_n
	);

	wire         clock_div_0_clk_neg_clk;                                        // clock_div_0:clk_neg -> [addr_delay_c_neg_0:pll_clock, addr_delay_c_neg_1:pll_clock, addr_delay_c_neg_2:pll_clock, addr_delay_c_neg_3:pll_clock, addr_delay_c_neg_4:pll_clock, dp_ram_a_neg:ram_clock, dp_ram_b_neg:ram_clock, dp_ram_c_neg:ram_clock, mc_data_delay_neg:div_clock, test_control_unit_0:pll_clock_neg]
	wire         clock_div_0_clk_pos_clk;                                        // clock_div_0:clk_pos -> [addr_delay_c_pos_0:pll_clock, addr_delay_c_pos_1:pll_clock, addr_delay_c_pos_2:pll_clock, addr_delay_c_pos_3:pll_clock, addr_delay_c_pos_4:pll_clock, dp_ram_a_pos:ram_clock, dp_ram_b_pos:ram_clock, dp_ram_c_pos:ram_clock, mc_data_delay_pos:div_clock, test_control_unit_0:pll_clock_pos]
	wire         pll_0_outclk0_clk;                                              // pll_0:outclk_0 -> [clock_div_0:clock, clocked_mux_a:clock, clocked_mux_b:clock, data_delay_a_0:pll_clock, data_delay_a_1:pll_clock, data_delay_b_0:pll_clock, data_delay_b_1:pll_clock, data_delay_neg_0:pll_clock, data_delay_neg_1:pll_clock, data_delay_pos_0:pll_clock, data_delay_pos_1:pll_clock, mc_data_delay_neg:pll_clock, mc_data_delay_pos:pll_clock, online_adder_0:clock]
	wire  [10:0] test_control_unit_0_read_a_neg_addr;                            // test_control_unit_0:r_addr_a_neg -> dp_ram_a_neg:addr_arith
	wire         test_control_unit_0_read_a_neg_we;                              // test_control_unit_0:we_read_a_neg -> dp_ram_a_neg:we_arith
	wire  [10:0] test_control_unit_0_read_a_pos_addr;                            // test_control_unit_0:r_addr_a_pos -> dp_ram_a_pos:addr_arith
	wire         test_control_unit_0_read_a_pos_we;                              // test_control_unit_0:we_read_a_pos -> dp_ram_a_pos:we_arith
	wire  [10:0] test_control_unit_0_read_b_neg_addr;                            // test_control_unit_0:r_addr_b_neg -> dp_ram_b_neg:addr_arith
	wire         test_control_unit_0_read_b_neg_we;                              // test_control_unit_0:we_read_b_neg -> dp_ram_b_neg:we_arith
	wire  [10:0] addr_delay_c_pos_0_addr_out_addr;                               // addr_delay_c_pos_0:addr_out -> addr_delay_c_pos_1:addr_in
	wire         addr_delay_c_pos_0_addr_out_we;                                 // addr_delay_c_pos_0:e_out -> addr_delay_c_pos_1:e_in
	wire  [10:0] addr_delay_c_neg_0_addr_out_addr;                               // addr_delay_c_neg_0:addr_out -> addr_delay_c_neg_1:addr_in
	wire         addr_delay_c_neg_0_addr_out_we;                                 // addr_delay_c_neg_0:e_out -> addr_delay_c_neg_1:e_in
	wire  [10:0] test_control_unit_0_write_neg_addr;                             // test_control_unit_0:w_addr_neg -> addr_delay_c_neg_0:addr_in
	wire         test_control_unit_0_write_neg_we;                               // test_control_unit_0:we_neg -> addr_delay_c_neg_0:e_in
	wire  [10:0] addr_delay_c_pos_4_addr_out_addr;                               // addr_delay_c_pos_4:addr_out -> dp_ram_c_pos:addr_arith
	wire         addr_delay_c_pos_4_addr_out_we;                                 // addr_delay_c_pos_4:e_out -> dp_ram_c_pos:we_arith
	wire  [10:0] addr_delay_c_neg_4_addr_out_addr;                               // addr_delay_c_neg_4:addr_out -> dp_ram_c_neg:addr_arith
	wire         addr_delay_c_neg_4_addr_out_we;                                 // addr_delay_c_neg_4:e_out -> dp_ram_c_neg:we_arith
	wire  [10:0] addr_delay_c_pos_1_addr_out_addr;                               // addr_delay_c_pos_1:addr_out -> addr_delay_c_pos_2:addr_in
	wire         addr_delay_c_pos_1_addr_out_we;                                 // addr_delay_c_pos_1:e_out -> addr_delay_c_pos_2:e_in
	wire  [10:0] addr_delay_c_neg_1_addr_out_addr;                               // addr_delay_c_neg_1:addr_out -> addr_delay_c_neg_2:addr_in
	wire         addr_delay_c_neg_1_addr_out_we;                                 // addr_delay_c_neg_1:e_out -> addr_delay_c_neg_2:e_in
	wire  [10:0] addr_delay_c_neg_2_addr_out_addr;                               // addr_delay_c_neg_2:addr_out -> addr_delay_c_neg_3:addr_in
	wire         addr_delay_c_neg_2_addr_out_we;                                 // addr_delay_c_neg_2:e_out -> addr_delay_c_neg_3:e_in
	wire  [10:0] addr_delay_c_pos_2_addr_out_addr;                               // addr_delay_c_pos_2:addr_out -> addr_delay_c_pos_3:addr_in
	wire         addr_delay_c_pos_2_addr_out_we;                                 // addr_delay_c_pos_2:e_out -> addr_delay_c_pos_3:e_in
	wire  [10:0] addr_delay_c_pos_3_addr_out_addr;                               // addr_delay_c_pos_3:addr_out -> addr_delay_c_pos_4:addr_in
	wire         addr_delay_c_pos_3_addr_out_we;                                 // addr_delay_c_pos_3:e_out -> addr_delay_c_pos_4:e_in
	wire  [10:0] addr_delay_c_neg_3_addr_out_addr;                               // addr_delay_c_neg_3:addr_out -> addr_delay_c_neg_4:addr_in
	wire         addr_delay_c_neg_3_addr_out_we;                                 // addr_delay_c_neg_3:e_out -> addr_delay_c_neg_4:e_in
	wire  [31:0] online_adder_0_c_out_data;                                      // online_adder_0:s_out -> arith_out_duplicate_0:data_in
	wire  [29:0] data_delay_a_1_data_out_data;                                   // data_delay_a_1:data_out -> online_adder_0:x_in
	wire  [29:0] data_delay_b_1_data_out_data;                                   // data_delay_b_1:data_out -> online_adder_0:y_in
	wire  [31:0] mc_data_delay_pos_data_out_data;                                // mc_data_delay_pos:data_out -> dp_ram_c_pos:data_arith
	wire  [31:0] mc_data_delay_neg_data_out_data;                                // mc_data_delay_neg:data_out -> dp_ram_c_neg:data_arith
	wire  [29:0] data_delay_a_0_data_out_data;                                   // data_delay_a_0:data_out -> data_delay_a_1:data_in
	wire  [29:0] data_delay_b_0_data_out_data;                                   // data_delay_b_0:data_out -> data_delay_b_1:data_in
	wire  [31:0] data_delay_pos_0_data_out_data;                                 // data_delay_pos_0:data_out -> data_delay_pos_1:data_in
	wire  [31:0] data_delay_pos_1_data_out_data;                                 // data_delay_pos_1:data_out -> mc_data_delay_pos:data_in
	wire  [31:0] data_delay_neg_0_data_out_data;                                 // data_delay_neg_0:data_out -> data_delay_neg_1:data_in
	wire  [31:0] data_delay_neg_1_data_out_data;                                 // data_delay_neg_1:data_out -> mc_data_delay_neg:data_in
	wire         pll_0_locked_export;                                            // pll_0:locked -> test_control_unit_0:pll_lock
	wire  [31:0] dp_ram_a_neg_q_arth_data;                                       // dp_ram_a_neg:q_arith -> clocked_mux_a:neg_in
	wire  [31:0] arith_out_duplicate_0_neg_out_data;                             // arith_out_duplicate_0:neg_out -> data_delay_neg_0:data_in
	wire  [31:0] dp_ram_b_pos_q_arth_data;                                       // dp_ram_b_pos:q_arith -> clocked_mux_b:pos_in
	wire  [31:0] arith_out_duplicate_0_pos_out_data;                             // arith_out_duplicate_0:pos_out -> data_delay_pos_0:data_in
	wire  [31:0] dp_ram_b_neg_q_arth_data;                                       // dp_ram_b_neg:q_arith -> clocked_mux_b:neg_in
	wire  [31:0] dp_ram_a_pos_q_arth_data;                                       // dp_ram_a_pos:q_arith -> clocked_mux_a:pos_in
	wire  [29:0] clocked_mux_a_q_out_data;                                       // clocked_mux_a:q_out -> data_delay_a_0:data_in
	wire  [29:0] clocked_mux_b_q_out_data;                                       // clocked_mux_b:q_out -> data_delay_b_0:data_in
	wire  [10:0] test_control_unit_0_read_b_pos_addr;                            // test_control_unit_0:r_addr_b_pos -> dp_ram_b_pos:addr_arith
	wire         test_control_unit_0_read_b_pos_we;                              // test_control_unit_0:we_read_b_pos -> dp_ram_b_pos:we_arith
	wire  [63:0] pll_0_reconfig_from_pll_reconfig_from_pll;                      // pll_0:reconfig_from_pll -> pll_reconfig_0:reconfig_from_pll
	wire  [63:0] pll_reconfig_0_reconfig_to_pll_reconfig_to_pll;                 // pll_reconfig_0:reconfig_to_pll -> pll_0:reconfig_to_pll
	wire  [10:0] test_control_unit_0_write_pos_addr;                             // test_control_unit_0:w_addr_pos -> addr_delay_c_pos_0:addr_in
	wire         test_control_unit_0_write_pos_we;                               // test_control_unit_0:we_pos -> addr_delay_c_pos_0:e_in
	wire   [1:0] hps_0_h2f_lw_axi_master_awburst;                                // hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	wire   [3:0] hps_0_h2f_lw_axi_master_arlen;                                  // hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	wire   [3:0] hps_0_h2f_lw_axi_master_wstrb;                                  // hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	wire         hps_0_h2f_lw_axi_master_wready;                                 // mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_rid;                                    // mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire         hps_0_h2f_lw_axi_master_rready;                                 // hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	wire   [3:0] hps_0_h2f_lw_axi_master_awlen;                                  // hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	wire  [11:0] hps_0_h2f_lw_axi_master_wid;                                    // hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	wire   [3:0] hps_0_h2f_lw_axi_master_arcache;                                // hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	wire         hps_0_h2f_lw_axi_master_wvalid;                                 // hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_0_h2f_lw_axi_master_araddr;                                 // hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	wire   [2:0] hps_0_h2f_lw_axi_master_arprot;                                 // hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	wire   [2:0] hps_0_h2f_lw_axi_master_awprot;                                 // hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	wire  [31:0] hps_0_h2f_lw_axi_master_wdata;                                  // hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	wire         hps_0_h2f_lw_axi_master_arvalid;                                // hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_0_h2f_lw_axi_master_awcache;                                // hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	wire  [11:0] hps_0_h2f_lw_axi_master_arid;                                   // hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	wire   [1:0] hps_0_h2f_lw_axi_master_arlock;                                 // hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	wire   [1:0] hps_0_h2f_lw_axi_master_awlock;                                 // hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	wire  [20:0] hps_0_h2f_lw_axi_master_awaddr;                                 // hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_0_h2f_lw_axi_master_bresp;                                  // mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire         hps_0_h2f_lw_axi_master_arready;                                // mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire  [31:0] hps_0_h2f_lw_axi_master_rdata;                                  // mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire         hps_0_h2f_lw_axi_master_awready;                                // mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [1:0] hps_0_h2f_lw_axi_master_arburst;                                // hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	wire   [2:0] hps_0_h2f_lw_axi_master_arsize;                                 // hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	wire         hps_0_h2f_lw_axi_master_bready;                                 // hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	wire         hps_0_h2f_lw_axi_master_rlast;                                  // mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire         hps_0_h2f_lw_axi_master_wlast;                                  // hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	wire   [1:0] hps_0_h2f_lw_axi_master_rresp;                                  // mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire  [11:0] hps_0_h2f_lw_axi_master_awid;                                   // hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	wire  [11:0] hps_0_h2f_lw_axi_master_bid;                                    // mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire         hps_0_h2f_lw_axi_master_bvalid;                                 // mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [2:0] hps_0_h2f_lw_axi_master_awsize;                                 // hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	wire         hps_0_h2f_lw_axi_master_awvalid;                                // hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	wire         hps_0_h2f_lw_axi_master_rvalid;                                 // mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire  [31:0] mm_interconnect_0_mm_bridge_0_s0_readdata;                      // mm_bridge_0:s0_readdata -> mm_interconnect_0:mm_bridge_0_s0_readdata
	wire         mm_interconnect_0_mm_bridge_0_s0_waitrequest;                   // mm_bridge_0:s0_waitrequest -> mm_interconnect_0:mm_bridge_0_s0_waitrequest
	wire         mm_interconnect_0_mm_bridge_0_s0_debugaccess;                   // mm_interconnect_0:mm_bridge_0_s0_debugaccess -> mm_bridge_0:s0_debugaccess
	wire  [10:0] mm_interconnect_0_mm_bridge_0_s0_address;                       // mm_interconnect_0:mm_bridge_0_s0_address -> mm_bridge_0:s0_address
	wire         mm_interconnect_0_mm_bridge_0_s0_read;                          // mm_interconnect_0:mm_bridge_0_s0_read -> mm_bridge_0:s0_read
	wire   [3:0] mm_interconnect_0_mm_bridge_0_s0_byteenable;                    // mm_interconnect_0:mm_bridge_0_s0_byteenable -> mm_bridge_0:s0_byteenable
	wire         mm_interconnect_0_mm_bridge_0_s0_readdatavalid;                 // mm_bridge_0:s0_readdatavalid -> mm_interconnect_0:mm_bridge_0_s0_readdatavalid
	wire         mm_interconnect_0_mm_bridge_0_s0_write;                         // mm_interconnect_0:mm_bridge_0_s0_write -> mm_bridge_0:s0_write
	wire  [31:0] mm_interconnect_0_mm_bridge_0_s0_writedata;                     // mm_interconnect_0:mm_bridge_0_s0_writedata -> mm_bridge_0:s0_writedata
	wire   [0:0] mm_interconnect_0_mm_bridge_0_s0_burstcount;                    // mm_interconnect_0:mm_bridge_0_s0_burstcount -> mm_bridge_0:s0_burstcount
	wire         mm_bridge_0_m0_waitrequest;                                     // mm_interconnect_1:mm_bridge_0_m0_waitrequest -> mm_bridge_0:m0_waitrequest
	wire  [31:0] mm_bridge_0_m0_readdata;                                        // mm_interconnect_1:mm_bridge_0_m0_readdata -> mm_bridge_0:m0_readdata
	wire         mm_bridge_0_m0_debugaccess;                                     // mm_bridge_0:m0_debugaccess -> mm_interconnect_1:mm_bridge_0_m0_debugaccess
	wire  [10:0] mm_bridge_0_m0_address;                                         // mm_bridge_0:m0_address -> mm_interconnect_1:mm_bridge_0_m0_address
	wire         mm_bridge_0_m0_read;                                            // mm_bridge_0:m0_read -> mm_interconnect_1:mm_bridge_0_m0_read
	wire   [3:0] mm_bridge_0_m0_byteenable;                                      // mm_bridge_0:m0_byteenable -> mm_interconnect_1:mm_bridge_0_m0_byteenable
	wire         mm_bridge_0_m0_readdatavalid;                                   // mm_interconnect_1:mm_bridge_0_m0_readdatavalid -> mm_bridge_0:m0_readdatavalid
	wire  [31:0] mm_bridge_0_m0_writedata;                                       // mm_bridge_0:m0_writedata -> mm_interconnect_1:mm_bridge_0_m0_writedata
	wire         mm_bridge_0_m0_write;                                           // mm_bridge_0:m0_write -> mm_interconnect_1:mm_bridge_0_m0_write
	wire   [0:0] mm_bridge_0_m0_burstcount;                                      // mm_bridge_0:m0_burstcount -> mm_interconnect_1:mm_bridge_0_m0_burstcount
	wire  [31:0] mm_interconnect_1_test_control_unit_0_avalon_slave_0_readdata;  // test_control_unit_0:readdata -> mm_interconnect_1:test_control_unit_0_avalon_slave_0_readdata
	wire   [2:0] mm_interconnect_1_test_control_unit_0_avalon_slave_0_address;   // mm_interconnect_1:test_control_unit_0_avalon_slave_0_address -> test_control_unit_0:address
	wire         mm_interconnect_1_test_control_unit_0_avalon_slave_0_read;      // mm_interconnect_1:test_control_unit_0_avalon_slave_0_read -> test_control_unit_0:read
	wire         mm_interconnect_1_test_control_unit_0_avalon_slave_0_write;     // mm_interconnect_1:test_control_unit_0_avalon_slave_0_write -> test_control_unit_0:write
	wire  [31:0] mm_interconnect_1_test_control_unit_0_avalon_slave_0_writedata; // mm_interconnect_1:test_control_unit_0_avalon_slave_0_writedata -> test_control_unit_0:writedata
	wire  [31:0] mm_interconnect_1_dp_ram_c_neg_avalon_slave_0_readdata;         // dp_ram_c_neg:readdata -> mm_interconnect_1:dp_ram_c_neg_avalon_slave_0_readdata
	wire   [4:0] mm_interconnect_1_dp_ram_c_neg_avalon_slave_0_address;          // mm_interconnect_1:dp_ram_c_neg_avalon_slave_0_address -> dp_ram_c_neg:address
	wire         mm_interconnect_1_dp_ram_c_neg_avalon_slave_0_read;             // mm_interconnect_1:dp_ram_c_neg_avalon_slave_0_read -> dp_ram_c_neg:read
	wire         mm_interconnect_1_dp_ram_c_neg_avalon_slave_0_write;            // mm_interconnect_1:dp_ram_c_neg_avalon_slave_0_write -> dp_ram_c_neg:write
	wire  [31:0] mm_interconnect_1_dp_ram_c_neg_avalon_slave_0_writedata;        // mm_interconnect_1:dp_ram_c_neg_avalon_slave_0_writedata -> dp_ram_c_neg:writedata
	wire  [31:0] mm_interconnect_1_dp_ram_c_pos_avalon_slave_0_readdata;         // dp_ram_c_pos:readdata -> mm_interconnect_1:dp_ram_c_pos_avalon_slave_0_readdata
	wire   [4:0] mm_interconnect_1_dp_ram_c_pos_avalon_slave_0_address;          // mm_interconnect_1:dp_ram_c_pos_avalon_slave_0_address -> dp_ram_c_pos:address
	wire         mm_interconnect_1_dp_ram_c_pos_avalon_slave_0_read;             // mm_interconnect_1:dp_ram_c_pos_avalon_slave_0_read -> dp_ram_c_pos:read
	wire         mm_interconnect_1_dp_ram_c_pos_avalon_slave_0_write;            // mm_interconnect_1:dp_ram_c_pos_avalon_slave_0_write -> dp_ram_c_pos:write
	wire  [31:0] mm_interconnect_1_dp_ram_c_pos_avalon_slave_0_writedata;        // mm_interconnect_1:dp_ram_c_pos_avalon_slave_0_writedata -> dp_ram_c_pos:writedata
	wire  [31:0] mm_interconnect_1_dp_ram_b_neg_avalon_slave_0_readdata;         // dp_ram_b_neg:readdata -> mm_interconnect_1:dp_ram_b_neg_avalon_slave_0_readdata
	wire   [4:0] mm_interconnect_1_dp_ram_b_neg_avalon_slave_0_address;          // mm_interconnect_1:dp_ram_b_neg_avalon_slave_0_address -> dp_ram_b_neg:address
	wire         mm_interconnect_1_dp_ram_b_neg_avalon_slave_0_read;             // mm_interconnect_1:dp_ram_b_neg_avalon_slave_0_read -> dp_ram_b_neg:read
	wire         mm_interconnect_1_dp_ram_b_neg_avalon_slave_0_write;            // mm_interconnect_1:dp_ram_b_neg_avalon_slave_0_write -> dp_ram_b_neg:write
	wire  [31:0] mm_interconnect_1_dp_ram_b_neg_avalon_slave_0_writedata;        // mm_interconnect_1:dp_ram_b_neg_avalon_slave_0_writedata -> dp_ram_b_neg:writedata
	wire  [31:0] mm_interconnect_1_dp_ram_b_pos_avalon_slave_0_readdata;         // dp_ram_b_pos:readdata -> mm_interconnect_1:dp_ram_b_pos_avalon_slave_0_readdata
	wire   [4:0] mm_interconnect_1_dp_ram_b_pos_avalon_slave_0_address;          // mm_interconnect_1:dp_ram_b_pos_avalon_slave_0_address -> dp_ram_b_pos:address
	wire         mm_interconnect_1_dp_ram_b_pos_avalon_slave_0_read;             // mm_interconnect_1:dp_ram_b_pos_avalon_slave_0_read -> dp_ram_b_pos:read
	wire         mm_interconnect_1_dp_ram_b_pos_avalon_slave_0_write;            // mm_interconnect_1:dp_ram_b_pos_avalon_slave_0_write -> dp_ram_b_pos:write
	wire  [31:0] mm_interconnect_1_dp_ram_b_pos_avalon_slave_0_writedata;        // mm_interconnect_1:dp_ram_b_pos_avalon_slave_0_writedata -> dp_ram_b_pos:writedata
	wire  [31:0] mm_interconnect_1_dp_ram_a_neg_avalon_slave_0_readdata;         // dp_ram_a_neg:readdata -> mm_interconnect_1:dp_ram_a_neg_avalon_slave_0_readdata
	wire   [4:0] mm_interconnect_1_dp_ram_a_neg_avalon_slave_0_address;          // mm_interconnect_1:dp_ram_a_neg_avalon_slave_0_address -> dp_ram_a_neg:address
	wire         mm_interconnect_1_dp_ram_a_neg_avalon_slave_0_read;             // mm_interconnect_1:dp_ram_a_neg_avalon_slave_0_read -> dp_ram_a_neg:read
	wire         mm_interconnect_1_dp_ram_a_neg_avalon_slave_0_write;            // mm_interconnect_1:dp_ram_a_neg_avalon_slave_0_write -> dp_ram_a_neg:write
	wire  [31:0] mm_interconnect_1_dp_ram_a_neg_avalon_slave_0_writedata;        // mm_interconnect_1:dp_ram_a_neg_avalon_slave_0_writedata -> dp_ram_a_neg:writedata
	wire  [31:0] mm_interconnect_1_dp_ram_a_pos_avalon_slave_0_readdata;         // dp_ram_a_pos:readdata -> mm_interconnect_1:dp_ram_a_pos_avalon_slave_0_readdata
	wire   [4:0] mm_interconnect_1_dp_ram_a_pos_avalon_slave_0_address;          // mm_interconnect_1:dp_ram_a_pos_avalon_slave_0_address -> dp_ram_a_pos:address
	wire         mm_interconnect_1_dp_ram_a_pos_avalon_slave_0_read;             // mm_interconnect_1:dp_ram_a_pos_avalon_slave_0_read -> dp_ram_a_pos:read
	wire         mm_interconnect_1_dp_ram_a_pos_avalon_slave_0_write;            // mm_interconnect_1:dp_ram_a_pos_avalon_slave_0_write -> dp_ram_a_pos:write
	wire  [31:0] mm_interconnect_1_dp_ram_a_pos_avalon_slave_0_writedata;        // mm_interconnect_1:dp_ram_a_pos_avalon_slave_0_writedata -> dp_ram_a_pos:writedata
	wire  [31:0] mm_interconnect_1_pll_reconfig_0_mgmt_avalon_slave_readdata;    // pll_reconfig_0:mgmt_readdata -> mm_interconnect_1:pll_reconfig_0_mgmt_avalon_slave_readdata
	wire         mm_interconnect_1_pll_reconfig_0_mgmt_avalon_slave_waitrequest; // pll_reconfig_0:mgmt_waitrequest -> mm_interconnect_1:pll_reconfig_0_mgmt_avalon_slave_waitrequest
	wire   [5:0] mm_interconnect_1_pll_reconfig_0_mgmt_avalon_slave_address;     // mm_interconnect_1:pll_reconfig_0_mgmt_avalon_slave_address -> pll_reconfig_0:mgmt_address
	wire         mm_interconnect_1_pll_reconfig_0_mgmt_avalon_slave_read;        // mm_interconnect_1:pll_reconfig_0_mgmt_avalon_slave_read -> pll_reconfig_0:mgmt_read
	wire         mm_interconnect_1_pll_reconfig_0_mgmt_avalon_slave_write;       // mm_interconnect_1:pll_reconfig_0_mgmt_avalon_slave_write -> pll_reconfig_0:mgmt_write
	wire  [31:0] mm_interconnect_1_pll_reconfig_0_mgmt_avalon_slave_writedata;   // mm_interconnect_1:pll_reconfig_0_mgmt_avalon_slave_writedata -> pll_reconfig_0:mgmt_writedata
	wire         rst_controller_reset_out_reset;                                 // rst_controller:reset_out -> [dp_ram_a_neg:resetn, dp_ram_a_pos:resetn, dp_ram_b_neg:resetn, dp_ram_b_pos:resetn, dp_ram_c_neg:resetn, dp_ram_c_pos:resetn, mm_bridge_0:reset, mm_interconnect_0:mm_bridge_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:mm_bridge_0_reset_reset_bridge_in_reset_reset, pll_reconfig_0:mgmt_reset, test_control_unit_0:resetn]
	wire         rst_controller_001_reset_out_reset;                             // rst_controller_001:reset_out -> mm_interconnect_0:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset

	addr_delay #(
		.ADDR_WIDTH (11)
	) addr_delay_c_neg_0 (
		.pll_clock (clock_div_0_clk_neg_clk),            //    clock.clk
		.addr_in   (test_control_unit_0_write_neg_addr), //  addr_in.addr
		.e_in      (test_control_unit_0_write_neg_we),   //         .we
		.addr_out  (addr_delay_c_neg_0_addr_out_addr),   // addr_out.addr
		.e_out     (addr_delay_c_neg_0_addr_out_we)      //         .we
	);

	addr_delay #(
		.ADDR_WIDTH (11)
	) addr_delay_c_neg_1 (
		.pll_clock (clock_div_0_clk_neg_clk),          //    clock.clk
		.addr_in   (addr_delay_c_neg_0_addr_out_addr), //  addr_in.addr
		.e_in      (addr_delay_c_neg_0_addr_out_we),   //         .we
		.addr_out  (addr_delay_c_neg_1_addr_out_addr), // addr_out.addr
		.e_out     (addr_delay_c_neg_1_addr_out_we)    //         .we
	);

	addr_delay #(
		.ADDR_WIDTH (11)
	) addr_delay_c_neg_2 (
		.pll_clock (clock_div_0_clk_neg_clk),          //    clock.clk
		.addr_in   (addr_delay_c_neg_1_addr_out_addr), //  addr_in.addr
		.e_in      (addr_delay_c_neg_1_addr_out_we),   //         .we
		.addr_out  (addr_delay_c_neg_2_addr_out_addr), // addr_out.addr
		.e_out     (addr_delay_c_neg_2_addr_out_we)    //         .we
	);

	addr_delay #(
		.ADDR_WIDTH (11)
	) addr_delay_c_neg_3 (
		.pll_clock (clock_div_0_clk_neg_clk),          //    clock.clk
		.addr_in   (addr_delay_c_neg_2_addr_out_addr), //  addr_in.addr
		.e_in      (addr_delay_c_neg_2_addr_out_we),   //         .we
		.addr_out  (addr_delay_c_neg_3_addr_out_addr), // addr_out.addr
		.e_out     (addr_delay_c_neg_3_addr_out_we)    //         .we
	);

	addr_delay #(
		.ADDR_WIDTH (11)
	) addr_delay_c_neg_4 (
		.pll_clock (clock_div_0_clk_neg_clk),          //    clock.clk
		.addr_in   (addr_delay_c_neg_3_addr_out_addr), //  addr_in.addr
		.e_in      (addr_delay_c_neg_3_addr_out_we),   //         .we
		.addr_out  (addr_delay_c_neg_4_addr_out_addr), // addr_out.addr
		.e_out     (addr_delay_c_neg_4_addr_out_we)    //         .we
	);

	addr_delay #(
		.ADDR_WIDTH (11)
	) addr_delay_c_pos_0 (
		.pll_clock (clock_div_0_clk_pos_clk),            //    clock.clk
		.addr_in   (test_control_unit_0_write_pos_addr), //  addr_in.addr
		.e_in      (test_control_unit_0_write_pos_we),   //         .we
		.addr_out  (addr_delay_c_pos_0_addr_out_addr),   // addr_out.addr
		.e_out     (addr_delay_c_pos_0_addr_out_we)      //         .we
	);

	addr_delay #(
		.ADDR_WIDTH (11)
	) addr_delay_c_pos_1 (
		.pll_clock (clock_div_0_clk_pos_clk),          //    clock.clk
		.addr_in   (addr_delay_c_pos_0_addr_out_addr), //  addr_in.addr
		.e_in      (addr_delay_c_pos_0_addr_out_we),   //         .we
		.addr_out  (addr_delay_c_pos_1_addr_out_addr), // addr_out.addr
		.e_out     (addr_delay_c_pos_1_addr_out_we)    //         .we
	);

	addr_delay #(
		.ADDR_WIDTH (11)
	) addr_delay_c_pos_2 (
		.pll_clock (clock_div_0_clk_pos_clk),          //    clock.clk
		.addr_in   (addr_delay_c_pos_1_addr_out_addr), //  addr_in.addr
		.e_in      (addr_delay_c_pos_1_addr_out_we),   //         .we
		.addr_out  (addr_delay_c_pos_2_addr_out_addr), // addr_out.addr
		.e_out     (addr_delay_c_pos_2_addr_out_we)    //         .we
	);

	addr_delay #(
		.ADDR_WIDTH (11)
	) addr_delay_c_pos_3 (
		.pll_clock (clock_div_0_clk_pos_clk),          //    clock.clk
		.addr_in   (addr_delay_c_pos_2_addr_out_addr), //  addr_in.addr
		.e_in      (addr_delay_c_pos_2_addr_out_we),   //         .we
		.addr_out  (addr_delay_c_pos_3_addr_out_addr), // addr_out.addr
		.e_out     (addr_delay_c_pos_3_addr_out_we)    //         .we
	);

	addr_delay #(
		.ADDR_WIDTH (11)
	) addr_delay_c_pos_4 (
		.pll_clock (clock_div_0_clk_pos_clk),          //    clock.clk
		.addr_in   (addr_delay_c_pos_3_addr_out_addr), //  addr_in.addr
		.e_in      (addr_delay_c_pos_3_addr_out_we),   //         .we
		.addr_out  (addr_delay_c_pos_4_addr_out_addr), // addr_out.addr
		.e_out     (addr_delay_c_pos_4_addr_out_we)    //         .we
	);

	arith_out_duplicate #(
		.IN_WIDTH  (32),
		.OUT_WIDTH (32)
	) arith_out_duplicate_0 (
		.neg_out (arith_out_duplicate_0_neg_out_data), // neg_out.data
		.pos_out (arith_out_duplicate_0_pos_out_data), // pos_out.data
		.data_in (online_adder_0_c_out_data)           // data_in.data
	);

	clock_div clock_div_0 (
		.clock   (pll_0_outclk0_clk),       // clock_sink.clk
		.clk_pos (clock_div_0_clk_pos_clk), //    clk_pos.clk
		.clk_neg (clock_div_0_clk_neg_clk)  //    clk_neg.clk
	);

	clocked_mux #(
		.IN_WIDTH  (32),
		.OUT_WIDTH (30),
		.INVERT    (1)
	) clocked_mux_a (
		.clock  (pll_0_outclk0_clk),        // clock_sink.clk
		.neg_in (dp_ram_a_neg_q_arth_data), //     neg_in.data
		.pos_in (dp_ram_a_pos_q_arth_data), //     pos_in.data
		.q_out  (clocked_mux_a_q_out_data)  //      q_out.data
	);

	clocked_mux #(
		.IN_WIDTH  (32),
		.OUT_WIDTH (30),
		.INVERT    (1)
	) clocked_mux_b (
		.clock  (pll_0_outclk0_clk),        // clock_sink.clk
		.neg_in (dp_ram_b_neg_q_arth_data), //     neg_in.data
		.pos_in (dp_ram_b_pos_q_arth_data), //     pos_in.data
		.q_out  (clocked_mux_b_q_out_data)  //      q_out.data
	);

	data_delay #(
		.WIDTH (30)
	) data_delay_a_0 (
		.pll_clock (pll_0_outclk0_clk),            //    clock.clk
		.data_in   (clocked_mux_a_q_out_data),     //  data_in.data
		.data_out  (data_delay_a_0_data_out_data)  // data_out.data
	);

	data_delay #(
		.WIDTH (30)
	) data_delay_a_1 (
		.pll_clock (pll_0_outclk0_clk),            //    clock.clk
		.data_in   (data_delay_a_0_data_out_data), //  data_in.data
		.data_out  (data_delay_a_1_data_out_data)  // data_out.data
	);

	data_delay #(
		.WIDTH (30)
	) data_delay_b_0 (
		.pll_clock (pll_0_outclk0_clk),            //    clock.clk
		.data_in   (clocked_mux_b_q_out_data),     //  data_in.data
		.data_out  (data_delay_b_0_data_out_data)  // data_out.data
	);

	data_delay #(
		.WIDTH (30)
	) data_delay_b_1 (
		.pll_clock (pll_0_outclk0_clk),            //    clock.clk
		.data_in   (data_delay_b_0_data_out_data), //  data_in.data
		.data_out  (data_delay_b_1_data_out_data)  // data_out.data
	);

	data_delay #(
		.WIDTH (32)
	) data_delay_neg_0 (
		.pll_clock (pll_0_outclk0_clk),                  //    clock.clk
		.data_in   (arith_out_duplicate_0_neg_out_data), //  data_in.data
		.data_out  (data_delay_neg_0_data_out_data)      // data_out.data
	);

	data_delay #(
		.WIDTH (32)
	) data_delay_neg_1 (
		.pll_clock (pll_0_outclk0_clk),              //    clock.clk
		.data_in   (data_delay_neg_0_data_out_data), //  data_in.data
		.data_out  (data_delay_neg_1_data_out_data)  // data_out.data
	);

	data_delay #(
		.WIDTH (32)
	) data_delay_pos_0 (
		.pll_clock (pll_0_outclk0_clk),                  //    clock.clk
		.data_in   (arith_out_duplicate_0_pos_out_data), //  data_in.data
		.data_out  (data_delay_pos_0_data_out_data)      // data_out.data
	);

	data_delay #(
		.WIDTH (32)
	) data_delay_pos_1 (
		.pll_clock (pll_0_outclk0_clk),              //    clock.clk
		.data_in   (data_delay_pos_0_data_out_data), //  data_in.data
		.data_out  (data_delay_pos_1_data_out_data)  // data_out.data
	);

	dpRam #(
		.ID         (3),
		.DATA_WIDTH (32),
		.ADDR_WIDTH (11)
	) dp_ram_a_neg (
		.resetn       (~rst_controller_reset_out_reset),                         //    clock_reset.reset_n
		.writedata    (mm_interconnect_1_dp_ram_a_neg_avalon_slave_0_writedata), // avalon_slave_0.writedata
		.readdata     (mm_interconnect_1_dp_ram_a_neg_avalon_slave_0_readdata),  //               .readdata
		.write        (mm_interconnect_1_dp_ram_a_neg_avalon_slave_0_write),     //               .write
		.read         (mm_interconnect_1_dp_ram_a_neg_avalon_slave_0_read),      //               .read
		.address      (mm_interconnect_1_dp_ram_a_neg_avalon_slave_0_address),   //               .address
		.avalon_clock (clk_clk),                                                 //     clock_sink.clk
		.ram_clock    (clock_div_0_clk_neg_clk),                                 //        pll_clk.clk
		.q_arith      (dp_ram_a_neg_q_arth_data),                                //         q_arth.data
		.data_arith   (),                                                        //      data_arth.data
		.addr_arith   (test_control_unit_0_read_a_neg_addr),                     //      addr_arth.addr
		.we_arith     (test_control_unit_0_read_a_neg_we)                        //               .we
	);

	dpRam #(
		.ID         (2),
		.DATA_WIDTH (32),
		.ADDR_WIDTH (11)
	) dp_ram_a_pos (
		.resetn       (~rst_controller_reset_out_reset),                         //    clock_reset.reset_n
		.writedata    (mm_interconnect_1_dp_ram_a_pos_avalon_slave_0_writedata), // avalon_slave_0.writedata
		.readdata     (mm_interconnect_1_dp_ram_a_pos_avalon_slave_0_readdata),  //               .readdata
		.write        (mm_interconnect_1_dp_ram_a_pos_avalon_slave_0_write),     //               .write
		.read         (mm_interconnect_1_dp_ram_a_pos_avalon_slave_0_read),      //               .read
		.address      (mm_interconnect_1_dp_ram_a_pos_avalon_slave_0_address),   //               .address
		.avalon_clock (clk_clk),                                                 //     clock_sink.clk
		.ram_clock    (clock_div_0_clk_pos_clk),                                 //        pll_clk.clk
		.q_arith      (dp_ram_a_pos_q_arth_data),                                //         q_arth.data
		.data_arith   (),                                                        //      data_arth.data
		.addr_arith   (test_control_unit_0_read_a_pos_addr),                     //      addr_arth.addr
		.we_arith     (test_control_unit_0_read_a_pos_we)                        //               .we
	);

	dpRam #(
		.ID         (5),
		.DATA_WIDTH (32),
		.ADDR_WIDTH (11)
	) dp_ram_b_neg (
		.resetn       (~rst_controller_reset_out_reset),                         //    clock_reset.reset_n
		.writedata    (mm_interconnect_1_dp_ram_b_neg_avalon_slave_0_writedata), // avalon_slave_0.writedata
		.readdata     (mm_interconnect_1_dp_ram_b_neg_avalon_slave_0_readdata),  //               .readdata
		.write        (mm_interconnect_1_dp_ram_b_neg_avalon_slave_0_write),     //               .write
		.read         (mm_interconnect_1_dp_ram_b_neg_avalon_slave_0_read),      //               .read
		.address      (mm_interconnect_1_dp_ram_b_neg_avalon_slave_0_address),   //               .address
		.avalon_clock (clk_clk),                                                 //     clock_sink.clk
		.ram_clock    (clock_div_0_clk_neg_clk),                                 //        pll_clk.clk
		.q_arith      (dp_ram_b_neg_q_arth_data),                                //         q_arth.data
		.data_arith   (),                                                        //      data_arth.data
		.addr_arith   (test_control_unit_0_read_b_neg_addr),                     //      addr_arth.addr
		.we_arith     (test_control_unit_0_read_b_neg_we)                        //               .we
	);

	dpRam #(
		.ID         (4),
		.DATA_WIDTH (32),
		.ADDR_WIDTH (11)
	) dp_ram_b_pos (
		.resetn       (~rst_controller_reset_out_reset),                         //    clock_reset.reset_n
		.writedata    (mm_interconnect_1_dp_ram_b_pos_avalon_slave_0_writedata), // avalon_slave_0.writedata
		.readdata     (mm_interconnect_1_dp_ram_b_pos_avalon_slave_0_readdata),  //               .readdata
		.write        (mm_interconnect_1_dp_ram_b_pos_avalon_slave_0_write),     //               .write
		.read         (mm_interconnect_1_dp_ram_b_pos_avalon_slave_0_read),      //               .read
		.address      (mm_interconnect_1_dp_ram_b_pos_avalon_slave_0_address),   //               .address
		.avalon_clock (clk_clk),                                                 //     clock_sink.clk
		.ram_clock    (clock_div_0_clk_pos_clk),                                 //        pll_clk.clk
		.q_arith      (dp_ram_b_pos_q_arth_data),                                //         q_arth.data
		.data_arith   (),                                                        //      data_arth.data
		.addr_arith   (test_control_unit_0_read_b_pos_addr),                     //      addr_arth.addr
		.we_arith     (test_control_unit_0_read_b_pos_we)                        //               .we
	);

	dpRam #(
		.ID         (7),
		.DATA_WIDTH (32),
		.ADDR_WIDTH (11)
	) dp_ram_c_neg (
		.resetn       (~rst_controller_reset_out_reset),                         //    clock_reset.reset_n
		.writedata    (mm_interconnect_1_dp_ram_c_neg_avalon_slave_0_writedata), // avalon_slave_0.writedata
		.readdata     (mm_interconnect_1_dp_ram_c_neg_avalon_slave_0_readdata),  //               .readdata
		.write        (mm_interconnect_1_dp_ram_c_neg_avalon_slave_0_write),     //               .write
		.read         (mm_interconnect_1_dp_ram_c_neg_avalon_slave_0_read),      //               .read
		.address      (mm_interconnect_1_dp_ram_c_neg_avalon_slave_0_address),   //               .address
		.avalon_clock (clk_clk),                                                 //     clock_sink.clk
		.ram_clock    (clock_div_0_clk_neg_clk),                                 //        pll_clk.clk
		.q_arith      (),                                                        //         q_arth.data
		.data_arith   (mc_data_delay_neg_data_out_data),                         //      data_arth.data
		.addr_arith   (addr_delay_c_neg_4_addr_out_addr),                        //      addr_arth.addr
		.we_arith     (addr_delay_c_neg_4_addr_out_we)                           //               .we
	);

	dpRam #(
		.ID         (6),
		.DATA_WIDTH (32),
		.ADDR_WIDTH (11)
	) dp_ram_c_pos (
		.resetn       (~rst_controller_reset_out_reset),                         //    clock_reset.reset_n
		.writedata    (mm_interconnect_1_dp_ram_c_pos_avalon_slave_0_writedata), // avalon_slave_0.writedata
		.readdata     (mm_interconnect_1_dp_ram_c_pos_avalon_slave_0_readdata),  //               .readdata
		.write        (mm_interconnect_1_dp_ram_c_pos_avalon_slave_0_write),     //               .write
		.read         (mm_interconnect_1_dp_ram_c_pos_avalon_slave_0_read),      //               .read
		.address      (mm_interconnect_1_dp_ram_c_pos_avalon_slave_0_address),   //               .address
		.avalon_clock (clk_clk),                                                 //     clock_sink.clk
		.ram_clock    (clock_div_0_clk_pos_clk),                                 //        pll_clk.clk
		.q_arith      (),                                                        //         q_arth.data
		.data_arith   (mc_data_delay_pos_data_out_data),                         //      data_arth.data
		.addr_arith   (addr_delay_c_pos_4_addr_out_addr),                        //      addr_arth.addr
		.we_arith     (addr_delay_c_pos_4_addr_out_we)                           //               .we
	);

	soc_system_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (0)
	) hps_0 (
		.mem_a                    (memory_mem_a),                          //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                         //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                         //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                       //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                        //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                       //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                      //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                      //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                       //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                    //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                         //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                        //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                      //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                        //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                         //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                      //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_0_hps_io_hps_io_emac1_inst_TX_CLK), //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_0_hps_io_hps_io_emac1_inst_TXD0),   //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_0_hps_io_hps_io_emac1_inst_TXD1),   //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_0_hps_io_hps_io_emac1_inst_TXD2),   //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_0_hps_io_hps_io_emac1_inst_TXD3),   //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_0_hps_io_hps_io_emac1_inst_RXD0),   //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_0_hps_io_hps_io_emac1_inst_MDIO),   //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_0_hps_io_hps_io_emac1_inst_MDC),    //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_0_hps_io_hps_io_emac1_inst_RX_CTL), //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_0_hps_io_hps_io_emac1_inst_TX_CTL), //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_0_hps_io_hps_io_emac1_inst_RX_CLK), //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_0_hps_io_hps_io_emac1_inst_RXD1),   //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_0_hps_io_hps_io_emac1_inst_RXD2),   //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_0_hps_io_hps_io_emac1_inst_RXD3),   //                  .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_0_hps_io_hps_io_qspi_inst_IO0),     //                  .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_0_hps_io_hps_io_qspi_inst_IO1),     //                  .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_0_hps_io_hps_io_qspi_inst_IO2),     //                  .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_0_hps_io_hps_io_qspi_inst_IO3),     //                  .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_0_hps_io_hps_io_qspi_inst_SS0),     //                  .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_0_hps_io_hps_io_qspi_inst_CLK),     //                  .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_0_hps_io_hps_io_sdio_inst_CMD),     //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_0_hps_io_hps_io_sdio_inst_D0),      //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_0_hps_io_hps_io_sdio_inst_D1),      //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_0_hps_io_hps_io_sdio_inst_CLK),     //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_0_hps_io_hps_io_sdio_inst_D2),      //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_0_hps_io_hps_io_sdio_inst_D3),      //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_0_hps_io_hps_io_usb1_inst_D0),      //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_0_hps_io_hps_io_usb1_inst_D1),      //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_0_hps_io_hps_io_usb1_inst_D2),      //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_0_hps_io_hps_io_usb1_inst_D3),      //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_0_hps_io_hps_io_usb1_inst_D4),      //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_0_hps_io_hps_io_usb1_inst_D5),      //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_0_hps_io_hps_io_usb1_inst_D6),      //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_0_hps_io_hps_io_usb1_inst_D7),      //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_0_hps_io_hps_io_usb1_inst_CLK),     //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_0_hps_io_hps_io_usb1_inst_STP),     //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_0_hps_io_hps_io_usb1_inst_DIR),     //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_0_hps_io_hps_io_usb1_inst_NXT),     //                  .hps_io_usb1_inst_NXT
		.hps_io_spim0_inst_CLK    (hps_0_hps_io_hps_io_spim0_inst_CLK),    //                  .hps_io_spim0_inst_CLK
		.hps_io_spim0_inst_MOSI   (hps_0_hps_io_hps_io_spim0_inst_MOSI),   //                  .hps_io_spim0_inst_MOSI
		.hps_io_spim0_inst_MISO   (hps_0_hps_io_hps_io_spim0_inst_MISO),   //                  .hps_io_spim0_inst_MISO
		.hps_io_spim0_inst_SS0    (hps_0_hps_io_hps_io_spim0_inst_SS0),    //                  .hps_io_spim0_inst_SS0
		.hps_io_uart0_inst_RX     (hps_0_hps_io_hps_io_uart0_inst_RX),     //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_0_hps_io_hps_io_uart0_inst_TX),     //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_0_hps_io_hps_io_i2c0_inst_SDA),     //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_0_hps_io_hps_io_i2c0_inst_SCL),     //                  .hps_io_i2c0_inst_SCL
		.hps_io_can0_inst_RX      (hps_0_hps_io_hps_io_can0_inst_RX),      //                  .hps_io_can0_inst_RX
		.hps_io_can0_inst_TX      (hps_0_hps_io_hps_io_can0_inst_TX),      //                  .hps_io_can0_inst_TX
		.hps_io_trace_inst_CLK    (hps_0_hps_io_hps_io_trace_inst_CLK),    //                  .hps_io_trace_inst_CLK
		.hps_io_trace_inst_D0     (hps_0_hps_io_hps_io_trace_inst_D0),     //                  .hps_io_trace_inst_D0
		.hps_io_trace_inst_D1     (hps_0_hps_io_hps_io_trace_inst_D1),     //                  .hps_io_trace_inst_D1
		.hps_io_trace_inst_D2     (hps_0_hps_io_hps_io_trace_inst_D2),     //                  .hps_io_trace_inst_D2
		.hps_io_trace_inst_D3     (hps_0_hps_io_hps_io_trace_inst_D3),     //                  .hps_io_trace_inst_D3
		.hps_io_trace_inst_D4     (hps_0_hps_io_hps_io_trace_inst_D4),     //                  .hps_io_trace_inst_D4
		.hps_io_trace_inst_D5     (hps_0_hps_io_hps_io_trace_inst_D5),     //                  .hps_io_trace_inst_D5
		.hps_io_trace_inst_D6     (hps_0_hps_io_hps_io_trace_inst_D6),     //                  .hps_io_trace_inst_D6
		.hps_io_trace_inst_D7     (hps_0_hps_io_hps_io_trace_inst_D7),     //                  .hps_io_trace_inst_D7
		.hps_io_gpio_inst_GPIO09  (hps_0_hps_io_hps_io_gpio_inst_GPIO09),  //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_0_hps_io_hps_io_gpio_inst_GPIO35),  //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO41  (hps_0_hps_io_hps_io_gpio_inst_GPIO41),  //                  .hps_io_gpio_inst_GPIO41
		.hps_io_gpio_inst_GPIO42  (hps_0_hps_io_hps_io_gpio_inst_GPIO42),  //                  .hps_io_gpio_inst_GPIO42
		.hps_io_gpio_inst_GPIO43  (hps_0_hps_io_hps_io_gpio_inst_GPIO43),  //                  .hps_io_gpio_inst_GPIO43
		.hps_io_gpio_inst_GPIO44  (hps_0_hps_io_hps_io_gpio_inst_GPIO44),  //                  .hps_io_gpio_inst_GPIO44
		.h2f_rst_n                (hps_0_h2f_reset_reset_n),               //         h2f_reset.reset_n
		.h2f_lw_axi_clk           (clk_clk),                               //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),          // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),        //                  .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),         //                  .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),        //                  .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst),       //                  .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),        //                  .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache),       //                  .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),        //                  .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid),       //                  .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready),       //                  .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),           //                  .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),         //                  .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),         //                  .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),         //                  .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),        //                  .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),        //                  .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),           //                  .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),         //                  .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),        //                  .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),        //                  .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),          //                  .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),        //                  .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),         //                  .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),        //                  .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst),       //                  .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),        //                  .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache),       //                  .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),        //                  .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid),       //                  .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready),       //                  .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),           //                  .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),         //                  .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),         //                  .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),         //                  .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),        //                  .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready)         //                  .rready
	);

	mc_data_delay #(
		.WIDTH  (32),
		.INVERT (0)
	) mc_data_delay_neg (
		.data_out  (mc_data_delay_neg_data_out_data), //  data_out.data
		.data_in   (data_delay_neg_1_data_out_data),  //   data_in.data
		.div_clock (clock_div_0_clk_neg_clk),         // div_clock.clk
		.pll_clock (pll_0_outclk0_clk)                // pll_clock.clk
	);

	mc_data_delay #(
		.WIDTH  (32),
		.INVERT (1)
	) mc_data_delay_pos (
		.data_out  (mc_data_delay_pos_data_out_data), //  data_out.data
		.data_in   (data_delay_pos_1_data_out_data),  //   data_in.data
		.div_clock (clock_div_0_clk_pos_clk),         // div_clock.clk
		.pll_clock (pll_0_outclk0_clk)                // pll_clock.clk
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (11),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_0 (
		.clk              (clk_clk),                                        //   clk.clk
		.reset            (rst_controller_reset_out_reset),                 // reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_bridge_0_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_bridge_0_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_bridge_0_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_bridge_0_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_mm_bridge_0_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_mm_bridge_0_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_mm_bridge_0_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_mm_bridge_0_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_mm_bridge_0_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_bridge_0_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mm_bridge_0_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (mm_bridge_0_m0_readdata),                        //      .readdata
		.m0_readdatavalid (mm_bridge_0_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (mm_bridge_0_m0_burstcount),                      //      .burstcount
		.m0_writedata     (mm_bridge_0_m0_writedata),                       //      .writedata
		.m0_address       (mm_bridge_0_m0_address),                         //      .address
		.m0_write         (mm_bridge_0_m0_write),                           //      .write
		.m0_read          (mm_bridge_0_m0_read),                            //      .read
		.m0_byteenable    (mm_bridge_0_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (mm_bridge_0_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                               // (terminated)
		.m0_response      (2'b00)                                           // (terminated)
	);

	rRp_add_clocked #(
		.RADIX (2),
		.WIDTH (15)
	) online_adder_0 (
		.x_in  (data_delay_a_1_data_out_data), //  a_in.data
		.y_in  (data_delay_b_1_data_out_data), //  b_in.data
		.s_out (online_adder_0_c_out_data),    // c_out.data
		.clock (pll_0_outclk0_clk)             // clock.clk
	);

	soc_system_pll_0 pll_0 (
		.refclk            (clk_clk),                                        //            refclk.clk
		.rst               (~reset_reset_n),                                 //             reset.reset
		.outclk_0          (pll_0_outclk0_clk),                              //           outclk0.clk
		.locked            (pll_0_locked_export),                            //            locked.export
		.reconfig_to_pll   (pll_reconfig_0_reconfig_to_pll_reconfig_to_pll), //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (pll_0_reconfig_from_pll_reconfig_from_pll)       // reconfig_from_pll.reconfig_from_pll
	);

	altera_pll_reconfig_top #(
		.device_family       ("Cyclone V"),
		.ENABLE_MIF          (0),
		.MIF_FILE_NAME       (""),
		.ENABLE_BYTEENABLE   (0),
		.BYTEENABLE_WIDTH    (4),
		.RECONFIG_ADDR_WIDTH (6),
		.RECONFIG_DATA_WIDTH (32),
		.reconf_width        (64),
		.WAIT_FOR_LOCK       (1)
	) pll_reconfig_0 (
		.mgmt_clk          (clk_clk),                                                        //          mgmt_clk.clk
		.mgmt_reset        (rst_controller_reset_out_reset),                                 //        mgmt_reset.reset
		.mgmt_waitrequest  (mm_interconnect_1_pll_reconfig_0_mgmt_avalon_slave_waitrequest), // mgmt_avalon_slave.waitrequest
		.mgmt_read         (mm_interconnect_1_pll_reconfig_0_mgmt_avalon_slave_read),        //                  .read
		.mgmt_write        (mm_interconnect_1_pll_reconfig_0_mgmt_avalon_slave_write),       //                  .write
		.mgmt_readdata     (mm_interconnect_1_pll_reconfig_0_mgmt_avalon_slave_readdata),    //                  .readdata
		.mgmt_address      (mm_interconnect_1_pll_reconfig_0_mgmt_avalon_slave_address),     //                  .address
		.mgmt_writedata    (mm_interconnect_1_pll_reconfig_0_mgmt_avalon_slave_writedata),   //                  .writedata
		.reconfig_to_pll   (pll_reconfig_0_reconfig_to_pll_reconfig_to_pll),                 //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (pll_0_reconfig_from_pll_reconfig_from_pll),                      // reconfig_from_pll.reconfig_from_pll
		.mgmt_byteenable   (4'b0000)                                                         //       (terminated)
	);

	testControlUnit #(
		.ID (8)
	) test_control_unit_0 (
		.writedata     (mm_interconnect_1_test_control_unit_0_avalon_slave_0_writedata), // avalon_slave_0.writedata
		.readdata      (mm_interconnect_1_test_control_unit_0_avalon_slave_0_readdata),  //               .readdata
		.write         (mm_interconnect_1_test_control_unit_0_avalon_slave_0_write),     //               .write
		.read          (mm_interconnect_1_test_control_unit_0_avalon_slave_0_read),      //               .read
		.address       (mm_interconnect_1_test_control_unit_0_avalon_slave_0_address),   //               .address
		.avalon_clock  (clk_clk),                                                        //     clock_sink.clk
		.resetn        (~rst_controller_reset_out_reset),                                //     reset_sink.reset_n
		.w_addr_pos    (test_control_unit_0_write_pos_addr),                             //      write_pos.addr
		.we_pos        (test_control_unit_0_write_pos_we),                               //               .we
		.w_addr_neg    (test_control_unit_0_write_neg_addr),                             //      write_neg.addr
		.we_neg        (test_control_unit_0_write_neg_we),                               //               .we
		.r_addr_a_pos  (test_control_unit_0_read_a_pos_addr),                            //     read_a_pos.addr
		.we_read_a_pos (test_control_unit_0_read_a_pos_we),                              //               .we
		.r_addr_a_neg  (test_control_unit_0_read_a_neg_addr),                            //     read_a_neg.addr
		.we_read_a_neg (test_control_unit_0_read_a_neg_we),                              //               .we
		.r_addr_b_pos  (test_control_unit_0_read_b_pos_addr),                            //     read_b_pos.addr
		.we_read_b_pos (test_control_unit_0_read_b_pos_we),                              //               .we
		.r_addr_b_neg  (test_control_unit_0_read_b_neg_addr),                            //     read_b_neg.addr
		.we_read_b_neg (test_control_unit_0_read_b_neg_we),                              //               .we
		.pll_clock_pos (clock_div_0_clk_pos_clk),                                        //  pll_clock_pos.clk
		.pll_clock_neg (clock_div_0_clk_neg_clk),                                        //  pll_clock_neg.clk
		.pll_lock      (pll_0_locked_export)                                             //       pll_lock.export
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                   //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                 //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                  //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                 //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                 //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                 //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                    //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                  //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                  //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                  //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                 //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                 //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                    //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                  //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                 //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                 //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                   //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                 //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                  //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                 //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                 //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                 //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                    //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                  //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                  //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                  //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                 //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                 //                                                              .rready
		.clk_0_clk_clk                                                       (clk_clk),                                        //                                                     clk_0_clk.clk
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),             // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_reset_reset_bridge_in_reset_reset                       (rst_controller_reset_out_reset),                 //                       mm_bridge_0_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_s0_address                                              (mm_interconnect_0_mm_bridge_0_s0_address),       //                                                mm_bridge_0_s0.address
		.mm_bridge_0_s0_write                                                (mm_interconnect_0_mm_bridge_0_s0_write),         //                                                              .write
		.mm_bridge_0_s0_read                                                 (mm_interconnect_0_mm_bridge_0_s0_read),          //                                                              .read
		.mm_bridge_0_s0_readdata                                             (mm_interconnect_0_mm_bridge_0_s0_readdata),      //                                                              .readdata
		.mm_bridge_0_s0_writedata                                            (mm_interconnect_0_mm_bridge_0_s0_writedata),     //                                                              .writedata
		.mm_bridge_0_s0_burstcount                                           (mm_interconnect_0_mm_bridge_0_s0_burstcount),    //                                                              .burstcount
		.mm_bridge_0_s0_byteenable                                           (mm_interconnect_0_mm_bridge_0_s0_byteenable),    //                                                              .byteenable
		.mm_bridge_0_s0_readdatavalid                                        (mm_interconnect_0_mm_bridge_0_s0_readdatavalid), //                                                              .readdatavalid
		.mm_bridge_0_s0_waitrequest                                          (mm_interconnect_0_mm_bridge_0_s0_waitrequest),   //                                                              .waitrequest
		.mm_bridge_0_s0_debugaccess                                          (mm_interconnect_0_mm_bridge_0_s0_debugaccess)    //                                                              .debugaccess
	);

	soc_system_mm_interconnect_1 mm_interconnect_1 (
		.clk_0_clk_clk                                 (clk_clk),                                                        //                               clk_0_clk.clk
		.mm_bridge_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                 // mm_bridge_0_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_m0_address                        (mm_bridge_0_m0_address),                                         //                          mm_bridge_0_m0.address
		.mm_bridge_0_m0_waitrequest                    (mm_bridge_0_m0_waitrequest),                                     //                                        .waitrequest
		.mm_bridge_0_m0_burstcount                     (mm_bridge_0_m0_burstcount),                                      //                                        .burstcount
		.mm_bridge_0_m0_byteenable                     (mm_bridge_0_m0_byteenable),                                      //                                        .byteenable
		.mm_bridge_0_m0_read                           (mm_bridge_0_m0_read),                                            //                                        .read
		.mm_bridge_0_m0_readdata                       (mm_bridge_0_m0_readdata),                                        //                                        .readdata
		.mm_bridge_0_m0_readdatavalid                  (mm_bridge_0_m0_readdatavalid),                                   //                                        .readdatavalid
		.mm_bridge_0_m0_write                          (mm_bridge_0_m0_write),                                           //                                        .write
		.mm_bridge_0_m0_writedata                      (mm_bridge_0_m0_writedata),                                       //                                        .writedata
		.mm_bridge_0_m0_debugaccess                    (mm_bridge_0_m0_debugaccess),                                     //                                        .debugaccess
		.dp_ram_a_neg_avalon_slave_0_address           (mm_interconnect_1_dp_ram_a_neg_avalon_slave_0_address),          //             dp_ram_a_neg_avalon_slave_0.address
		.dp_ram_a_neg_avalon_slave_0_write             (mm_interconnect_1_dp_ram_a_neg_avalon_slave_0_write),            //                                        .write
		.dp_ram_a_neg_avalon_slave_0_read              (mm_interconnect_1_dp_ram_a_neg_avalon_slave_0_read),             //                                        .read
		.dp_ram_a_neg_avalon_slave_0_readdata          (mm_interconnect_1_dp_ram_a_neg_avalon_slave_0_readdata),         //                                        .readdata
		.dp_ram_a_neg_avalon_slave_0_writedata         (mm_interconnect_1_dp_ram_a_neg_avalon_slave_0_writedata),        //                                        .writedata
		.dp_ram_a_pos_avalon_slave_0_address           (mm_interconnect_1_dp_ram_a_pos_avalon_slave_0_address),          //             dp_ram_a_pos_avalon_slave_0.address
		.dp_ram_a_pos_avalon_slave_0_write             (mm_interconnect_1_dp_ram_a_pos_avalon_slave_0_write),            //                                        .write
		.dp_ram_a_pos_avalon_slave_0_read              (mm_interconnect_1_dp_ram_a_pos_avalon_slave_0_read),             //                                        .read
		.dp_ram_a_pos_avalon_slave_0_readdata          (mm_interconnect_1_dp_ram_a_pos_avalon_slave_0_readdata),         //                                        .readdata
		.dp_ram_a_pos_avalon_slave_0_writedata         (mm_interconnect_1_dp_ram_a_pos_avalon_slave_0_writedata),        //                                        .writedata
		.dp_ram_b_neg_avalon_slave_0_address           (mm_interconnect_1_dp_ram_b_neg_avalon_slave_0_address),          //             dp_ram_b_neg_avalon_slave_0.address
		.dp_ram_b_neg_avalon_slave_0_write             (mm_interconnect_1_dp_ram_b_neg_avalon_slave_0_write),            //                                        .write
		.dp_ram_b_neg_avalon_slave_0_read              (mm_interconnect_1_dp_ram_b_neg_avalon_slave_0_read),             //                                        .read
		.dp_ram_b_neg_avalon_slave_0_readdata          (mm_interconnect_1_dp_ram_b_neg_avalon_slave_0_readdata),         //                                        .readdata
		.dp_ram_b_neg_avalon_slave_0_writedata         (mm_interconnect_1_dp_ram_b_neg_avalon_slave_0_writedata),        //                                        .writedata
		.dp_ram_b_pos_avalon_slave_0_address           (mm_interconnect_1_dp_ram_b_pos_avalon_slave_0_address),          //             dp_ram_b_pos_avalon_slave_0.address
		.dp_ram_b_pos_avalon_slave_0_write             (mm_interconnect_1_dp_ram_b_pos_avalon_slave_0_write),            //                                        .write
		.dp_ram_b_pos_avalon_slave_0_read              (mm_interconnect_1_dp_ram_b_pos_avalon_slave_0_read),             //                                        .read
		.dp_ram_b_pos_avalon_slave_0_readdata          (mm_interconnect_1_dp_ram_b_pos_avalon_slave_0_readdata),         //                                        .readdata
		.dp_ram_b_pos_avalon_slave_0_writedata         (mm_interconnect_1_dp_ram_b_pos_avalon_slave_0_writedata),        //                                        .writedata
		.dp_ram_c_neg_avalon_slave_0_address           (mm_interconnect_1_dp_ram_c_neg_avalon_slave_0_address),          //             dp_ram_c_neg_avalon_slave_0.address
		.dp_ram_c_neg_avalon_slave_0_write             (mm_interconnect_1_dp_ram_c_neg_avalon_slave_0_write),            //                                        .write
		.dp_ram_c_neg_avalon_slave_0_read              (mm_interconnect_1_dp_ram_c_neg_avalon_slave_0_read),             //                                        .read
		.dp_ram_c_neg_avalon_slave_0_readdata          (mm_interconnect_1_dp_ram_c_neg_avalon_slave_0_readdata),         //                                        .readdata
		.dp_ram_c_neg_avalon_slave_0_writedata         (mm_interconnect_1_dp_ram_c_neg_avalon_slave_0_writedata),        //                                        .writedata
		.dp_ram_c_pos_avalon_slave_0_address           (mm_interconnect_1_dp_ram_c_pos_avalon_slave_0_address),          //             dp_ram_c_pos_avalon_slave_0.address
		.dp_ram_c_pos_avalon_slave_0_write             (mm_interconnect_1_dp_ram_c_pos_avalon_slave_0_write),            //                                        .write
		.dp_ram_c_pos_avalon_slave_0_read              (mm_interconnect_1_dp_ram_c_pos_avalon_slave_0_read),             //                                        .read
		.dp_ram_c_pos_avalon_slave_0_readdata          (mm_interconnect_1_dp_ram_c_pos_avalon_slave_0_readdata),         //                                        .readdata
		.dp_ram_c_pos_avalon_slave_0_writedata         (mm_interconnect_1_dp_ram_c_pos_avalon_slave_0_writedata),        //                                        .writedata
		.pll_reconfig_0_mgmt_avalon_slave_address      (mm_interconnect_1_pll_reconfig_0_mgmt_avalon_slave_address),     //        pll_reconfig_0_mgmt_avalon_slave.address
		.pll_reconfig_0_mgmt_avalon_slave_write        (mm_interconnect_1_pll_reconfig_0_mgmt_avalon_slave_write),       //                                        .write
		.pll_reconfig_0_mgmt_avalon_slave_read         (mm_interconnect_1_pll_reconfig_0_mgmt_avalon_slave_read),        //                                        .read
		.pll_reconfig_0_mgmt_avalon_slave_readdata     (mm_interconnect_1_pll_reconfig_0_mgmt_avalon_slave_readdata),    //                                        .readdata
		.pll_reconfig_0_mgmt_avalon_slave_writedata    (mm_interconnect_1_pll_reconfig_0_mgmt_avalon_slave_writedata),   //                                        .writedata
		.pll_reconfig_0_mgmt_avalon_slave_waitrequest  (mm_interconnect_1_pll_reconfig_0_mgmt_avalon_slave_waitrequest), //                                        .waitrequest
		.test_control_unit_0_avalon_slave_0_address    (mm_interconnect_1_test_control_unit_0_avalon_slave_0_address),   //      test_control_unit_0_avalon_slave_0.address
		.test_control_unit_0_avalon_slave_0_write      (mm_interconnect_1_test_control_unit_0_avalon_slave_0_write),     //                                        .write
		.test_control_unit_0_avalon_slave_0_read       (mm_interconnect_1_test_control_unit_0_avalon_slave_0_read),      //                                        .read
		.test_control_unit_0_avalon_slave_0_readdata   (mm_interconnect_1_test_control_unit_0_avalon_slave_0_readdata),  //                                        .readdata
		.test_control_unit_0_avalon_slave_0_writedata  (mm_interconnect_1_test_control_unit_0_avalon_slave_0_writedata)  //                                        .writedata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
