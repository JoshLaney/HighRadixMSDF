module add_tester(
	avalon clk, pll_clk, clk_pos, clk_neg,
	
)